`timescale 1ns/1ps

module and_gate_tb;
    reg a, b;
    wire y;

    and_gate uut (
        .a(a),
        .b(b),
        .y(y)
    );

    initial begin
        // This creates a file for viewing waveforms
        $dumpfile("dump.vcd");
        $dumpvars(0, and_gate_tb);

        $display("A B | Y");
        $display("---------");
        
        a = 0; b = 0; #10; $display("%b %b | %b", a, b, y);
        a = 0; b = 1; #10; $display("%b %b | %b", a, b, y);
        a = 1; b = 0; #10; $display("%b %b | %b", a, b, y);
        a = 1; b = 1; #10; $display("%b %b | %b", a, b, y);
        
        $finish;
    end
endmodule
